library IEEE;
use IEEE.std_logic_1164.all;

entity TopFrame
	port();
end;

architecture  struct of  TopFrame is
begin

end;
